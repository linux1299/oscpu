`include "defines.v"

module axi_master_if # (
    parameter RW_DATA_WIDTH     = 64,
    parameter RW_ADDR_WIDTH     = 64,
    parameter AXI_DATA_WIDTH    = 64,
    parameter AXI_ADDR_WIDTH    = 64,
    parameter AXI_ID_WIDTH      = 4,
    parameter AXI_USER_WIDTH    = 1
)(
    input                               clk,
    input                               rst_n,

    // user port
    input                               rw_id_i,
    input                               rw_cen_i,
    input                               rw_wen_i,
    input  [RW_ADDR_WIDTH-1:0]          rw_addr_i,
    input  [2:0]                        rw_size_i,
    input  [RW_DATA_WIDTH-1:0]          rw_wdata_i,
    input  [7:0]                        rw_wmask_i,
    output                              rw_ready_o,
    output [RW_DATA_WIDTH-1:0]          rw_rdata_o,
    output [1:0]                        rw_resp_o,

    //------------AXI port-------------------------
    // write address channel
    output [AXI_ID_WIDTH-1:0]           axi_aw_id_o,
    output [AXI_ADDR_WIDTH-1:0]         axi_aw_addr_o,
    output [7:0]                        axi_aw_len_o,
    output [2:0]                        axi_aw_size_o,
    output [1:0]                        axi_aw_burst_o,
    output                              axi_aw_lock_o,
    output [3:0]                        axi_aw_cache_o,
    output [2:0]                        axi_aw_prot_o,
    output [3:0]                        axi_aw_qos_o,
    output [3:0]                        axi_aw_region_o,
    output [AXI_USER_WIDTH-1:0]         axi_aw_user_o,
    output                              axi_aw_valid_o,
    input                               axi_aw_ready_i,

    // write data channel
    input                               axi_w_ready_i,
    output                              axi_w_valid_o,
    output [AXI_DATA_WIDTH-1:0]         axi_w_data_o,
    output [AXI_DATA_WIDTH/8-1:0]       axi_w_strb_o,
    output                              axi_w_last_o,
    output [AXI_USER_WIDTH-1:0]         axi_w_user_o,

    // write response channel
    output                              axi_b_ready_o,
    input                               axi_b_valid_i,
    input  [1:0]                        axi_b_resp_i,
    input  [AXI_ID_WIDTH-1:0]           axi_b_id_i,
    input  [AXI_USER_WIDTH-1:0]         axi_b_user_i,

    // read address channel
    input                               axi_ar_ready_i,
    output                              axi_ar_valid_o,
    output [AXI_ADDR_WIDTH-1:0]         axi_ar_addr_o,
    output [2:0]                        axi_ar_prot_o,
    output [AXI_ID_WIDTH-1:0]           axi_ar_id_o,
    output [AXI_USER_WIDTH-1:0]         axi_ar_user_o,
    output [7:0]                        axi_ar_len_o,
    output [2:0]                        axi_ar_size_o,
    output [1:0]                        axi_ar_burst_o,
    output                              axi_ar_lock_o,
    output [3:0]                        axi_ar_cache_o,
    output [3:0]                        axi_ar_qos_o,
    output [3:0]                        axi_ar_region_o,

    // read data channel
    output                              axi_r_ready_o,
    input                               axi_r_valid_i,
    input  [1:0]                        axi_r_resp_i,
    input  [AXI_DATA_WIDTH-1:0]         axi_r_data_i,
    input                               axi_r_last_i,
    input  [AXI_ID_WIDTH-1:0]           axi_r_id_i,
    input  [AXI_USER_WIDTH-1:0]         axi_r_user_i
);

wire w_trans    = rw_wen_i;
wire r_trans    = ~rw_wen_i;
wire w_valid    = rw_cen_i & w_trans;
wire r_valid    = rw_cen_i & r_trans;

// handshake
wire aw_hs      = axi_aw_ready_i & axi_aw_valid_o;
wire w_hs       = axi_w_ready_i  & axi_w_valid_o;
wire b_hs       = axi_b_ready_o  & axi_b_valid_i;
wire ar_hs      = axi_ar_ready_i & axi_ar_valid_o;
wire r_hs       = axi_r_ready_o  & axi_r_valid_i;

wire w_done     = w_hs & axi_w_last_o;
wire r_done     = r_hs & axi_r_last_i;
wire trans_done = w_trans ? b_hs : r_done;


// ------------------State Machine------------------
localparam [2:0] W_STATE_IDLE  = 3'b000;
localparam [2:0] W_STATE_ADDR  = 3'b001;
localparam [2:0] W_STATE_WRITE = 3'b010;
localparam [2:0] W_STATE_RESP  = 3'b011;
localparam [2:0] W_STATE_DONE  = 3'b100;

localparam [1:0] R_STATE_IDLE  = 2'b00;
localparam [1:0] R_STATE_ADDR  = 2'b01;
localparam [1:0] R_STATE_READ  = 2'b10;
localparam [1:0] R_STATE_DONE  = 2'b11;

reg [2:0] w_state;
reg [1:0] r_state;

wire w_state_idle  = w_state == W_STATE_IDLE;
wire w_state_addr  = w_state == W_STATE_ADDR;
wire w_state_write = w_state == W_STATE_WRITE;
wire w_state_resp  = w_state == W_STATE_RESP;
wire w_state_done  = w_state == W_STATE_DONE;

wire r_state_idle  = r_state == R_STATE_IDLE;
wire r_state_addr  = r_state == R_STATE_ADDR;
wire r_state_read  = r_state == R_STATE_READ;
wire r_state_done  = r_state == R_STATE_DONE;

// ------------ Wirte State Machine --------------
always @(posedge clk) begin
    if (~rst_n) begin
        w_state <= W_STATE_IDLE;
    end
    else begin
        if (w_valid) begin
            case (w_state)
                W_STATE_IDLE:               w_state <= W_STATE_ADDR;
                W_STATE_ADDR:  if (aw_hs)   w_state <= W_STATE_WRITE;
                W_STATE_WRITE: if (w_done)  w_state <= W_STATE_RESP;
                W_STATE_RESP:  if (b_hs)    w_state <= W_STATE_DONE;
                W_STATE_DONE:               w_state <= W_STATE_IDLE;
            endcase
        end
    end
end

// ----------------- Read State Machine ----------------
always @(posedge clk) begin
    if (~rst_n) begin
        r_state <= R_STATE_IDLE;
    end
    else begin
        if (r_valid) begin
            case (r_state)
                R_STATE_IDLE:               r_state <= R_STATE_ADDR;
                R_STATE_ADDR: if (ar_hs)    r_state <= R_STATE_READ;
                R_STATE_READ: if (r_done)   r_state <= R_STATE_DONE;
                R_STATE_DONE:               r_state <= R_STATE_IDLE;
                default:;
            endcase
        end
    end
end




// ------------------Write Transaction------------------
// Write address channel signals
wire [AXI_ID_WIDTH-1:0]   axi_id   = {AXI_ID_WIDTH{1'b0}};
wire [AXI_USER_WIDTH-1:0] axi_user = {AXI_USER_WIDTH{1'b0}};
assign axi_aw_id_o      = axi_id;
assign axi_aw_addr_o    = rw_addr_i;
assign axi_aw_len_o     = 8'd0;
assign axi_aw_size_o    = rw_size_i;
assign axi_aw_burst_o   = `AXI_BURST_TYPE_INCR;
assign axi_aw_lock_o    = 1'b0;
assign axi_aw_cache_o   = `AXI_ARCACHE_NORMAL_NON_CACHEABLE_NON_BUFFERABLE;
assign axi_aw_prot_o    = `AXI_PROT_UNPRIVILEGED_ACCESS;
assign axi_aw_qos_o     = 4'h0;
assign axi_aw_region_o  = 4'h0;
assign axi_aw_user_o    = axi_user;
assign axi_aw_valid_o   = w_state_addr;

// Write data channel signals
assign axi_w_valid_o    = w_state_write;
assign axi_w_data_o     = rw_wdata_i;
assign axi_w_strb_o     = rw_wmask_i;
assign axi_w_last_o     = w_state_write;
assign axi_w_user_o     = axi_user;

// Write resp channel signals
assign axi_b_ready_o    = w_state_resp;


// ------------------Read Transaction------------------
// Read address channel signals
assign axi_ar_valid_o   = r_state_addr;
assign axi_ar_addr_o    = rw_addr_i;
assign axi_ar_prot_o    = `AXI_PROT_UNPRIVILEGED_ACCESS;
assign axi_ar_id_o      = axi_id;
assign axi_ar_user_o    = axi_user;
assign axi_ar_len_o     = 8'd0;
assign axi_ar_size_o    = rw_size_i;
assign axi_ar_burst_o   = `AXI_BURST_TYPE_INCR;
assign axi_ar_lock_o    = 1'b0;
assign axi_ar_cache_o   = `AXI_ARCACHE_NORMAL_NON_CACHEABLE_NON_BUFFERABLE;
assign axi_ar_qos_o     = 4'h0;

// Read data channel signals
assign axi_r_ready_o    = r_state_read;


// ------------------User Ports------------------
assign rw_rdata_o = axi_r_data_i;

reg  rw_ready;
always @(posedge clk) begin
    if (~rst_n) begin
        rw_ready <= 0;
    end
    else if (trans_done) begin
        rw_ready <= 1;
    end
    else begin
        rw_ready <= 0;
    end
end
assign rw_ready_o = rw_ready;

reg [1:0] rw_resp;
wire      rw_resp_next = w_trans ? axi_b_resp_i : axi_r_resp_i;
always @(posedge clk) begin
    if (~rst_n) begin
        rw_resp <= 0;
    end
    else if (trans_done) begin
        rw_resp <= rw_resp_next;
    end
    else begin
        rw_resp <= 0;
    end
end
assign rw_resp_o = rw_resp;


endmodule